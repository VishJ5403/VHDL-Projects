library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;

entity test is
end entity test;

architecture arc of test is
	constant ilen : integer := 16;		--length of instruction in bits
	
	component DUT is
		port (I: in std_logic_vector(ilen-1 downto 0); Iw,clk,iclk: in std_logic);
	end component DUT;

	signal I : std_logic_vector(ilen-1 downto 0);
	signal Iw : std_logic := '1';					--Instruction write
	signal clk: std_logic := '0';
	signal iclk: std_logic := '0';

	function to_string(x: string) return string is
		variable ret_val : string(1 to x'length);
		alias lx : string(1 to x'length) is x;
	begin
		ret_val := lx;
		return ret_val;
	end to_string;

	function to_std_logic_vector(x: bit_vector) return std_logic_vector is
		variable ret_val : std_logic_vector(1 to x'length);
		alias lx : bit_vector(1 to x'length) is x;
	begin
		for i in 1 to x'length loop
			if (lx(i)='1') then
				ret_val(i) := '1';
			else
				ret_val(i) := '0';
			end if;
		end loop;
		return ret_val;
	end to_std_logic_vector;

	function to_bit_vector(x: std_logic_vector) return bit_vector is
		variable ret_val : bit_vector(1 to x'length);
		alias lx : std_logic_vector(1 to x'length) is x;
	begin
		for i in 1 to x'length loop
			if (lx(i)='1') then
				ret_val(i) := '1';
			else
				ret_val(i) := '0';
			end if;
		end loop;
		return ret_val;
	end to_bit_vector;

begin
	process
		File infile : text open read_mode is "PROGRAM.txt";
		variable I_var : bit_vector(ilen-1 downto 0);
		variable input_line : line;
		variable line_count : integer := 0;
	begin
		while not endfile(infile) loop
			line_count := line_count + 1;
			readline (infile,input_line);
			read (input_line, I_var);
			I <= to_std_logic_vector(I_var);
			wait for 5 ns;
		end loop;
		Iw <= '0';
		wait;
	end process;
	
	iclock : process
	begin
		wait for 5 ns;
		iclk <= not iclk;
	end process;

	clock : process
	begin
		if (Iw = '1') then
			wait for 163840 ns;
		end if;
		wait for 5 ns;
		clk <= not clk;
	end process;

	DUT0 : DUT port map (I,Iw,clk,iclk);
end arc;

