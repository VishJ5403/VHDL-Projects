library ieee;
use ieee.std_logic_1164.all;

package memory_dm is
	component mem_dm is
		port (I,A,Din: in std_logic_vector(15 downto 0); Iw,r,w,clk,iclk: in std_logic; Dout: out std_logic_vector(15 downto 0));
	end component mem_dm;
end package memory_dm;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mem_dm is
	port (I,A,Din: in std_logic_vector(15 downto 0); Iw,r,w,clk,iclk:in std_logic; Dout: out std_logic_vector(15 downto 0));
end entity mem_dm;

architecture arc of mem_dm is
	type mem_array is array (0 to 65535) of std_logic_vector(15 downto 0);
	signal m: mem_array;
begin
--	process (I,Iw,iclk)
--		variable l: integer := 0;
--	begin
--		if (Iw='1') then
--			m(l) <= I;
--			l := l+1;
--		end if;
--	end process;
	process (A,Din,r,w,iclk,clk)
		variable l: integer := 0;
	begin
			if (Iw='1') then
				m(l) <= I;
				l := l+1;
			else
				if (r='1' AND w='0') then
				--address = (to_integer(unsigned(A)));
					Dout(15 downto 0) <= m(to_integer(unsigned(A)));		--big endian
				--Dout(7 downto 0) <= m((2*to_integer(unsigned(A)))+1);
				elsif(r='0' AND w='1') then
					if(clk'event and clk='0') then
					--address = to_integer(unsigned(A));
						m(to_integer(unsigned(A))) <= Din(15 downto 0);		--big endian
					--m((2*to_integer(unsigned(A)))+1) <= Din(7 downto 0);
					end if;
				end if;
			end if;
	end process;
end arc;
